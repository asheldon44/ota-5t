.save @n.x1.xm1a.nsg13_lv_nmos[ids] 
.save @n.x1.xm1a.nsg13_lv_nmos[vth]
.save @n.x1.xm1a.nsg13_lv_nmos[gm] 
.save @n.x1.xm1a.nsg13_lv_nmos[gmb] 
.save @n.x1.xm1a.nsg13_lv_nmos[gds] 
.save @n.x1.xm1a.nsg13_lv_nmos[cgg]
.save @n.x1.xm1a.nsg13_lv_nmos[cgs]
.save @n.x1.xm1a.nsg13_lv_nmos[cgd]
.save @n.x1.xm1a.nsg13_lv_nmos[cgb]
.save @n.x1.xm1a.nsg13_lv_nmos[cdd]
.save @n.x1.xm1a.nsg13_lv_nmos[css]
.save @n.x1.xm1a.nsg13_lv_nmos[cgsol]
.save @n.x1.xm1a.nsg13_lv_nmos[cgdol]
.save @n.x1.xm1a.nsg13_lv_nmos[cjs]
.save @n.x1.xm1a.nsg13_lv_nmos[cjd]
.save @n.x1.xm1a.nsg13_lv_nmos[vsat]
.save @n.x1.xm1b.nsg13_lv_nmos[ids]
.save @n.x1.xm1b.nsg13_lv_nmos[vth]
.save @n.x1.xm1b.nsg13_lv_nmos[gm]
.save @n.x1.xm1b.nsg13_lv_nmos[gmb]
.save @n.x1.xm1b.nsg13_lv_nmos[gds]
.save @n.x1.xm1b.nsg13_lv_nmos[cgg]
.save @n.x1.xm1b.nsg13_lv_nmos[cgs]
.save @n.x1.xm1b.nsg13_lv_nmos[cgd]
.save @n.x1.xm1b.nsg13_lv_nmos[cgb]
.save @n.x1.xm1b.nsg13_lv_nmos[cdd]
.save @n.x1.xm1b.nsg13_lv_nmos[css]
.save @n.x1.xm1b.nsg13_lv_nmos[cgsol]
.save @n.x1.xm1b.nsg13_lv_nmos[cgdol]
.save @n.x1.xm1b.nsg13_lv_nmos[cjs]
.save @n.x1.xm1b.nsg13_lv_nmos[cjd]
.save @n.x1.xm1b.nsg13_lv_nmos[vsat]
.save @n.x1.xm2a.nsg13_lv_pmos[ids]
.save @n.x1.xm2a.nsg13_lv_pmos[vth]
.save @n.x1.xm2a.nsg13_lv_pmos[gm]
.save @n.x1.xm2a.nsg13_lv_pmos[gmb]
.save @n.x1.xm2a.nsg13_lv_pmos[gds]
.save @n.x1.xm2a.nsg13_lv_pmos[cgg]
.save @n.x1.xm2a.nsg13_lv_pmos[cgs]
.save @n.x1.xm2a.nsg13_lv_pmos[cgd]
.save @n.x1.xm2a.nsg13_lv_pmos[cgb]
.save @n.x1.xm2a.nsg13_lv_pmos[cdd]
.save @n.x1.xm2a.nsg13_lv_pmos[css]
.save @n.x1.xm2a.nsg13_lv_pmos[cgsol]
.save @n.x1.xm2a.nsg13_lv_pmos[cgdol]
.save @n.x1.xm2a.nsg13_lv_pmos[cjs]
.save @n.x1.xm2a.nsg13_lv_pmos[cjd]
.save @n.x1.xm2a.nsg13_lv_pmos[vsat]
.save @n.x1.xm2b.nsg13_lv_pmos[ids]
.save @n.x1.xm2b.nsg13_lv_pmos[vth]
.save @n.x1.xm2b.nsg13_lv_pmos[gm]
.save @n.x1.xm2b.nsg13_lv_pmos[gmb]
.save @n.x1.xm2b.nsg13_lv_pmos[gds]
.save @n.x1.xm2b.nsg13_lv_pmos[cgg]
.save @n.x1.xm2b.nsg13_lv_pmos[cgs]
.save @n.x1.xm2b.nsg13_lv_pmos[cgd]
.save @n.x1.xm2b.nsg13_lv_pmos[cgb]
.save @n.x1.xm2b.nsg13_lv_pmos[cdd]
.save @n.x1.xm2b.nsg13_lv_pmos[css]
.save @n.x1.xm2b.nsg13_lv_pmos[cgsol]
.save @n.x1.xm2b.nsg13_lv_pmos[cgdol]
.save @n.x1.xm2b.nsg13_lv_pmos[cjs]
.save @n.x1.xm2b.nsg13_lv_pmos[cjd]
.save @n.x1.xm2b.nsg13_lv_pmos[vsat]
