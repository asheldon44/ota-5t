** sch_path: /foss/designs/ota_5t/ota-5t.sch
**.subckt ota-5t Vp Vn Vout VDD VSS Ib
*.iopin VDD
*.ipin Vn
*.opin Vout
*.ipin Vp
*.iopin VSS
*.ipin Ib
Xm1a vd Vn vs VSS sg13_lv_nmos w=10u l=4u ng=1 m=4
Xm2b vint vd VDD VDD sg13_lv_pmos w=2u l=2u ng=1 m=1
Xm2a vd vd VDD VDD sg13_lv_pmos w=2u l=2u ng=1 m=1
Xm3a vs Ib VSS VSS sg13_lv_nmos w=1u l=1u ng=1 m=2
Xm1b vint Vp vs VSS sg13_lv_nmos w=10u l=4u ng=1 m=4
Xm3ref Ib Ib VSS VSS sg13_lv_nmos w=1u l=1u ng=1 m=2
Xm3b vint2 Ib VSS VSS sg13_lv_nmos w=1u l=1u ng=1 m=2
Xm2c vint2 vint VDD VDD sg13_lv_pmos w=4u l=1u ng=1 m=1
Xm2d VDD vint2 Vout Vout sg13_lv_nmos w=1u l=1u ng=1 m=64
Xm3c Vout Ib VSS VSS sg13_lv_nmos w=1u l=1u ng=1 m=8
**.ends
.end
