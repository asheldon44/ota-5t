** sch_path: /foss/pdks/sg13g2/libs.tech/xschem/sg13g2_tests/dc_lv_nmos.sch
**.subckt dc_lv_nmos
Vgs net1 GND 0.75
Vds net3 GND 1.5
Vd net3 net2 0
.save i(vd)
XM1 net2 net1 GND GND sg13_lv_nmos w=12.7u l=0.13u ng=2 m=1
**** begin user architecture code
 .lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt



.param temp=27
.control
save all
op
*reset
dc Vds 0 3 0.01 Vgs 0. 0.9 0.1
write dc_lv_nmos.raw
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
