** sch_path: /foss/designs/ota_5t/tb_ota_5t_hier.sch
**.subckt tb_ota_5t_hier
Vin vin GND dc 0.6 ac 1
Vdd VDD GND 1.2
.save i(vdd)
C1 vout GND 1p m=1
x1 vin vout vout VDD GND net1 ota-5t
I1 VDD net1 10u
**** begin user architecture code
 .lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt



.param temp=27
.include /foss/designs/ota_5t/tb_ota_5t_save.spice
.control
	save all
	op
	write tb_ota_5t_hier.raw
	dc Vin 0 1.2 0.05
	plot v(vout) v(vin)
	plot v(vout)-v(vin)
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/ota_5t/ota-5t.sym # of pins=6
** sym_path: /foss/designs/ota_5t/ota-5t.sym
** sch_path: /foss/designs/ota_5t/ota-5t.sch
.subckt ota-5t Vp Vn Vout VDD VSS Ib
*.iopin VDD
*.ipin Vp
*.opin Vout
*.ipin Vn
*.iopin VSS
*.ipin Ib
Xm1a vd Vp vs VSS sg13_lv_nmos w=10u l=4u ng=1 m=4
Xm2b Vout vd VDD VDD sg13_lv_pmos w=2u l=2u ng=1 m=2
Xm2a vd vd VDD VDD sg13_lv_pmos w=2u l=2u ng=1 m=2
Xm3a vs Ib VSS VSS sg13_lv_nmos w=10u l=10u ng=1 m=2
Xm1b Vout Vn vs VSS sg13_lv_nmos w=10u l=4u ng=1 m=4
Xm3b Ib Ib VSS VSS sg13_lv_nmos w=10u l=10u ng=1 m=2
.ends

.GLOBAL GND
.end
