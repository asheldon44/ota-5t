** sch_path: /foss/designs/ota_5t/ota-5t_tb.sch
**.subckt ota-5t_tb
x1 vin net1 vout VDD GND net2 ota-5t
x999 net1 vout sub_x999
.subckt sub_x999 a b
Ii 0 x DC 0 AC 0
Vi x a DC 0 AC 1
Vnodebuffer b x 0
.ends loopgainprobe

.func tian_loop() {1/(1-1/(2*(ac1.I(v.X999.Vi)*ac2.V(X999.x)-ac1.V(X999.x)*ac2.I(v.X999.Vi))+ac1.V(X999.x)+ac2.I(v.X999.Vi)))}

C1 vout GND 1p m=1
Vin vin GND 0.6
Vsup VDD GND 1.2
I0 VDD net2 5u
**** begin user architecture code


 .lib /foss/pdks/sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt




.param temp=27
.include /foss/designs/ota_5t/tb_ota_5t_save.spice
.control
        save all
        op
        write ota-5t_tb.raw
        dc Vin 0 1.2 0.05
        plot v(vout) v(vin)
        plot v(vout)-v(vin)
        alter Vin 0.6
        ac dec 100 0.01 100e9
        alter i.X999.ii acmag=1
        alter v.X999.vi acmag=1
        ac dec 100 0.01 100e9
        let tian_signal = tian_loop()
        plot db(tian_signal)
        let dbsignal = db(tian_signal)
        meas ac zerogainfreq when dbsignal=0
        plot 180*cph(tian_signal)/pi
        let tphase = 180*cph(tian_signal)/pi
        meas ac phaseatzerogain find tphase at=zerogainfreq
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /foss/designs/ota_5t/ota-5t.sym # of pins=6
** sym_path: /foss/designs/ota_5t/ota-5t.sym
** sch_path: /foss/designs/ota_5t/ota-5t.sch
.subckt ota-5t Vp Vn Vout VDD VSS Ib
*.iopin VDD
*.ipin Vp
*.opin Vout
*.ipin Vn
*.iopin VSS
*.ipin Ib
Xm1a vd Vp vs VSS sg13_lv_nmos w=10u l=4u ng=1 m=4
Xm2b Vout vd VDD VDD sg13_lv_pmos w=2u l=1u ng=1 m=1
Xm2a vd vd VDD VDD sg13_lv_pmos w=2u l=1u ng=1 m=1
Xm3a vs Ib VSS VSS sg13_lv_nmos w=1u l=1u ng=1 m=2
Xm1b Vout Vn vs VSS sg13_lv_nmos w=10u l=4u ng=1 m=4
Xm3b Ib Ib VSS VSS sg13_lv_nmos w=1u l=1u ng=1 m=2
.ends

.GLOBAL GND
.end
